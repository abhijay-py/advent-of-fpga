module top (
    input logic clk,
    input logic rst_n,
    input logic serial_direction, // 1 = right, 0 = left
    input logic [15:0] serial_distance, // how many clicks to turn the dial
    output logic [15:0] password
)


endmodule